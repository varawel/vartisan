module vartisan

pub fn create_new()
{
	println("new")
}
